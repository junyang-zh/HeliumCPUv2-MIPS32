// forward.v: handles the pipeline forwarding

module forward (
    input wire idex_rs_reg_read, idex_rt_reg_read,
    input wire idex_rs_addr, idex_rt_addr,
    input wire exmem_reg_write,
    input wire exmem_write_dst
);
    
endmodule