// writeback.v

`include "defines.v"

module writeback (
    
);
    
endmodule